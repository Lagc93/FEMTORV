module uart_tx #(
    parameter CLK_FREQ = 27000000,
    parameter BAUD_RATE = 115200
)(
    input  wire clk,
    input  wire rst_n,
    input  wire tx_start,
    input  wire [7:0] tx_data,
    output reg  tx,
    output reg  tx_busy
);

    localparam DIV_CNT = CLK_FREQ / BAUD_RATE;

    reg [15:0] div_cnt;
    reg [3:0]  bit_cnt;
    reg [9:0]  tx_shift;

    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            tx       <= 1'b1;
            tx_busy  <= 0;
            div_cnt  <= 0;
            bit_cnt  <= 0;
            tx_shift <= 10'b1111111111;
        end else begin
            if (tx_start && !tx_busy) begin
                tx_shift <= {1'b1, tx_data, 1'b0}; // stop + data + start
                tx_busy  <= 1;
                bit_cnt  <= 0;
                div_cnt  <= 0;
            end else if (tx_busy) begin
                if (div_cnt == DIV_CNT-1) begin
                    div_cnt <= 0;
                    tx      <= tx_shift[bit_cnt];
                    bit_cnt <= bit_cnt + 1;
                    if (bit_cnt == 9) begin
                        tx_busy <= 0;
                    end
                end else begin
                    div_cnt <= div_cnt + 1;
                end
            end
        end
    end
endmodule
